module tb_regfile();

reg clk;
reg reset;  
