module tb_regfile();

reg clk;
reg reset;  

// TODO: Setup clock

// TOOD: Test regfile

    // TODO: Use monitor statement to display all register values

    // TODO: Test reset

    // TODO: Test writing to a single register

    // TODO: Test writing to multiple registers
        // TODO: Make sure not all registers get the bus value
    
    // TODO: Test output value aligns with desired register value
